module FreqDivHL(output reg sel0, sel1);
always @(*)begin
sel0 = 0;
sel1 = 1;
end
endmodule